//
// Author: <AUTHORNAME> (<AUTHOREMAIL>)
// Committer: <COMMITTERNAME>
//
// Creation Date:  Sat Apr 8 21:13:17 GMT+2 2017
// Module Name:    J1ScNexys4DDR - Behavioral
// Project Name:   J1Sc - A simple J1 implementation in Scala using Spinal HDL
//
// Hash: <COMMITHASH>
// Date: <AUTHORDATE>
//

module J1ScNexys4DDR (reset,
		      clk100Mhz, 
		      extInt,
		      leds,   
		      pmodA,
		      rx,    
		      tx);

 // Input ports
 input reset;
 input clk100Mhz;
 input [0:0] extInt;
 input rx;

 // Output ports
 output [15:0] leds;
 output tx;

 // Bidirectional port
 inout [7:0] pmodA;

 // Internal wiring 
 wire [7:0] pmodA_read;
 wire [7:0] pmodA_write;
 wire [7:0] pmodA_writeEnable;

 // Instantiate the J1SoC core generated by Spinal
 J1SoC core (.reset              (reset),
             .clk100Mhz          (clk100Mhz),
             .extInt             (extInt),
             .leds               (leds),
             .pmodA_read         (pmodA_read),
             .pmodA_write        (pmodA_write),
             .pmodA_writeEnable  (pmodA_writeEnable),
             .rx                 (rx),
             .tx                 (tx));

  // Connect the pmodA read port
  pmodA_read = pmodA;

  // Generate the write port and equip it with tristate functionality
  genvar i;
  generate 
     for (i = 0; i < 8; i = i + 1) begin
	assign pmodA[i] = pmodA_writeEnable[i] ? pmodA_write[i] : 1'bZ;
  end

endmodule // End of J1ScNexys4DDR
