//
// Author: Steffen Reith (steffen.reith@hs-rm.de)
//
// Creation Date:  Sat May 6 16:32:24 GMT+2 2017 
// Module Name:    Board_Nexys4 - Behavioral
// Project Name:   J1Sc - A simple J1 implementation in Scala using Spinal HDL
//
//

module Board_Nexys4 (reset,
		     clk100Mhz, 
 		     extInt,
		     leds,
                     rgbLeds,
                     segments_a,
                     segments_b,
                     segments_c,
                     segments_d,
                     segments_e,
                     segments_f,		     
                     segments_g,
                     dot,
                     selector,   
           	     pmodA,
		     sSwitches,
		     pButtons,
		     rx,    
		     tx);
		                
 // Input ports
 input reset;
 input clk100Mhz;
 input [0:0] extInt;
 input [15:0] sSwitches;  
 input [4:0] pButtons;  
 input rx;

 // Output ports
 output [15:0] leds;
 output tx;
 output segments_a;  
 output segments_b;  
 output segments_c; 
 output segments_d;  
 output segments_e;  
 output segments_f;  
 output segments_g;  
 output dot; 
 output [7:0] selector;

 // Bidirectional port
 inout [7:0] pmodA;

 // Clock generation
 wire boardClk;
 wire boardClkLocked;

 // Internal wiring 
 wire [7:0] pmodA_read;
 wire [7:0] pmodA_write;
 wire [7:0] pmodA_writeEnable;

 // Instantiate a PLL/MMCM (makes a 80Mhz clock)
 PLL makeClk (.clkIn    (clk100Mhz),
              .clkOut   (boardClk),
              .isLocked (boardClkLocked));

 // Instantiate the J1SoC core generated by Spinal
 J1SoC core (.reset              (reset),
             .boardClk           (boardClk),
             .boardClkLocked     (boardClkLocked),
             .extInt             (extInt),
             .leds               (leds),
             .rgbLeds            (rgbLeds),
             .segments_a         (segments_a),
             .segments_b         (segments_b),
             .segments_c         (segments_c),
             .segments_d         (segments_d),
             .segments_e         (segments_e),
             .segments_f         (segments_f),
             .segments_g         (segments_g),
	     .dot                (dot),
	     .selector           (selector),
             .pmodA_read         (pmodA_read),
             .pmodA_write        (pmodA_write),
             .pmodA_writeEnable  (pmodA_writeEnable),
	     .sSwitches          (sSwitches),
	     .pButtons           (pButtons),
             .rx                 (rx),
             .tx                 (tx));

  // Connect the pmodA read port
  assign pmodA_read = pmodA;

  // Generate the write port and equip it with tristate functionality
  genvar i;
  generate
     for (i = 0; i < 8; i = i + 1) begin
	   assign pmodA[i] = pmodA_writeEnable[i] ? pmodA_write[i] : 1'bZ;
     end
  endgenerate
  
endmodule

